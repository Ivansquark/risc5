module rv_alu( 
	input clkin,
	output clkout
);

assign clkout = clkin;



endmodule 