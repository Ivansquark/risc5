module decoder



endmodule;
